//Gabriel Altman
//ECEN2350 Digital Logic
//April, 2018

module Project_2_TOP
(
	MAX10_CLK1_50,
	MAX10_CLK2_50,
	LEDR,
	HEX0,
	HEX1,
	HEX2,
	HEX3,
	HEX4,
	HEX5,
	KEY,
	SW
);


input			MAX10_CLK1_50;						//50Mhz system clock 1
input			MAX10_CLK2_50;						//50Mhz system clock 2
input	[1:0]	KEY;									//Push-Buttons
input	[9:0]	SW;									//Switches

output	[9:0]	LEDR;								//LED's (Surface mounted) 
output	[7:0]	HEX0;								//Seven segment display 0
output	[7:0]	HEX1;								//Seven segment display 0
output	[7:0]	HEX2;								//Seven segment display 0
output	[7:0]	HEX3;								//Seven segment display 0
output	[7:0]	HEX4;								//Seven segment display 0
output	[7:0]	HEX5;								//Seven segment display 0

wire [1:0]ENABLE;									//Enable boolean
wire [1:0]RESET;									//Reset boolean
wire [3:0]BCD0;									//BCD 0
wire [3:0]BCD1;									//BCD 1
wire [3:0]BCD2;									//BCD 2
wire [3:0]BCD3;									//BCD 3
wire [9:0]divided_Clock;						//the 2kHz clock signal
wire [9:0]Slow_Clock;							//The 1Hz clock signal
wire [7:0]LFSR_Value;							//The random number generated by the LSFR
wire [1:0]downCount_Complete;					//boolean indicating the down_Counter has completed its count
wire [7:0]count;									//the value returned by the down_Counter showing the current value
wire [1:0]counter_Enable;						//boolean to enable the counter
wire [1:0]down_CounterEnable;					//boolean to enable the down_Counter


assign ENABLE[0] = SW[0];
assign RESET[0] = !KEY[0];

//Instantiates an instance of SevenSegment.v
//This is the decoder which translates BCD values into binary values that light the correct segments in the 7-segment display
BCD_decoder decoder_INST1(BCD0[3:0], BCD1[3:0], BCD2[3:0], BCD3[3:0], HEX0[6:0], HEX1[6:0], HEX2[6:0], HEX3[6:0]);

//Instantiates an instance of BCD_counter.v
//This code generates the values which generate numbers 1-9 for the seven-segment displays
BCD_counter BCD_Count_INST1(divided_Clock, RESET, ENABLE, BCD3, BCD2, BCD1, BCD0);

//Instantiates an instance of Clock_divider
//This clock divides the native 50MHz clock by 25,000 to yield a 2kHz clock
clock_Divider clk_Div_INST1(MAX10_CLK1_50, divided_Clock);

//Instantiates an instance of Slow_Clock
//This clock divides the native 50MHz clock by 50,000,000 to yield a 1Hz clock
Slow_Clock Slow_Clock_INST1(MAX10_CLK1_50, Slow_Clock);

//Instantiates an instance  of LFSR 
//Generates pseudo random numbers to set the delay between pressing the start button, and the start of the timer/start indicator light
LFSR LFSR_INST1(Slow_Clock, LFSR_Value);

//instantiates an instance of down_Counter
//down_Counter down_Counter_INST1(Slow_Clock, LFSR_Value, RESET, ENABLE, count, downCount_Complete);
down_Counter down_Counter_INST1(Slow_Clock, 8'b00000011, RESET, ENABLE, count, downCount_Complete);

assign HEX0[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display
assign HEX1[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display
assign HEX2[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display
assign HEX3[7] = 1'b0;						//Turns ON the decimal point for the 7-segment display
assign HEX4[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display
assign HEX5[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display

assign HEX4 = 8'b11111111;					//Blanks digit 4 of the 7-segment display
assign HEX5 = 8'b11111111;					//Blanks digit 5 of the 7-segment display

assign LEDR[9] = !KEY[0];					//TEMPORARY indicator for the reset switch
assign LEDR[8] = downCount_Complete;	//TEMPORARY indicator for the downCount_Complete boolean 1=count complete
//assign LEDR[7:0] = LFSR_Value[7:0];	//TEMPORARY indicator to verify the operation of the LSFR_Value module (Pseudo-Random number generator)
assign LEDR[7:0] = count[7:0];			//TEMPORARY indicator to verify the operation of the down_Counter module

endmodule
