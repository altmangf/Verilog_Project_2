//Gabriel Altman
//ECEN2350 Digital Logic
//April, 2018

module Project_2_TOP
(
	MAX10_CLK1_50,
	MAX10_CLK2_50,
	LEDR,
	HEX0,
	HEX1,
	HEX2,
	HEX3,
	HEX4,
	HEX5,
	KEY,
	SW
);


input			MAX10_CLK1_50;						//50Mhz system clock 1
input			MAX10_CLK2_50;						//50Mhz system clock 2
input	[1:0]	KEY;									//Push-Buttons
input	[9:0]	SW;									//Switches

output	[9:0]	LEDR;								//LED's (Surface mounted) 
output	[7:0]	HEX0;								//Seven segment display 0
output	[7:0]	HEX1;								//Seven segment display 0
output	[7:0]	HEX2;								//Seven segment display 0
output	[7:0]	HEX3;								//Seven segment display 0
output	[7:0]	HEX4;								//Seven segment display 0
output	[7:0]	HEX5;								//Seven segment display 0

reg [1:0]ENABLE;									//Enable boolean
wire [1:0]RESET;									//Reset boolean
wire [3:0]BCD0;									//BCD 0
wire [3:0]BCD1;									//BCD 1
wire [3:0]BCD2;									//BCD 2
wire [3:0]BCD3;									//BCD 3
wire [9:0]divided_Clock;						//the 2kHz clock signal
wire [9:0]Slow_Clock;							//The 1Hz clock signal
wire [7:0]LFSR_Value;							//The random number generated by the LSFR
wire [1:0]downCount_Complete;					//boolean indicating the down_Counter has completed its count
wire [7:0]count;									//the value returned by the down_Counter showing the current value
reg [1:0]counter_Enable;						//boolean to enable the counter
reg [1:0]downCounter_Enable;					//boolean to enable the down_Counter
reg [15:0]highScore;								//High score
reg [15:0]currentScore;							//current score
reg [2:0]A;											//Current state of Finite State Machine
reg downCount_Boolean;							//count complete=1  count running=0
reg downCount_Value;								//The LFSR value assigned to the down counter
 
//assign ENABLE[0] = SW[0];
assign RESET[0] = !KEY[0];					//Toggles the RESET boolean
assign HEX0[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display
assign HEX1[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display
assign HEX2[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display
assign HEX3[7] = 1'b0;						//Turns ON the decimal point for the 7-segment display
assign HEX4[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display
assign HEX5[7] = 1'b1;						//Turns OFF the decimal point for the 7-segment display
assign HEX4 = 8'b11111111;					//Blanks digit 4 of the 7-segment display
assign HEX5 = 8'b11111111;					//Blanks digit 5 of the 7-segment display
assign LEDR[9] = !KEY[0];					//indicator for the reset switch
assign LEDR[8] = downCount_Complete;	//indicator for the downCount_Complete boolean 1=count complete
assign LEDR[7] = downCount_Complete;	//indicator for the downCount_Complete boolean 1=count complete
assign LEDR[6] = downCount_Complete;	//indicator for the downCount_Complete boolean 1=count complete
assign LEDR[5] = downCount_Complete;	//indicator for the downCount_Complete boolean 1=count complete
assign LEDR[4] = downCount_Complete;	//indicator for the downCount_Complete boolean 1=count complete
//assign LEDR[7:0] = LFSR_Value[7:0];	//TEMPORARY indicator to verify the operation of the LSFR_Value module (Pseudo-Random number generator)
//assign LEDR[7:0] = count[7:0];			//TEMPORARY indicator to verify the operation of the down_Counter module
//assign downCount_Boolean = downCount_Complete;
assign LEDR[2:0] = A[2:0];					//TEMPORARY indicator to show current state of FSM 


/*always@(KEY[0])
begin
	if(KEY[0]==0)
		ENABLE = !ENABLE;
	if(KEY[1]==0)
		highScore = 0;
		A=2'b00;
		counter_Enable = 0;
		downCounter_Enable = 0;
		downCount_Boolean = 0;
end
*/



always@(A, KEY[1], KEY[0], SW[9], downCount_Boolean, downCount_Complete)
begin
	if(KEY[0]==0)begin
		highScore <= 0;
		A<=3'b000;
		counter_Enable <= 0;
		downCounter_Enable <= 0;
		downCount_Boolean <= 0;
		A <= 0;
		end
	//if(A == 3'b000 && SW[9] ==1'b0 && KEY[1] == 1'b1)begin
		//A <= 3'b001;
		//counter_Enable <= 0;
		//downCounter_Enable <=0;
		//downCount_Complete <=0;
		//display High Score
		//end
	if(A == 3'b000 && SW[9] ==1'b0 && KEY[1] == 1'b0)begin
		A <= 3'b001;
		counter_Enable <= 0;
		downCounter_Enable <=0;
		//downCount_Complete <=0;
		//display High Score
		end
	else if(A == 3'b000 && SW[9] == 1'b1 && KEY[1] == 1'b1)begin
		A <= 3'b111;
		counter_Enable <= 0;
		downCounter_Enable <=0;
		//downCount_Complete <=0;
		//Display "Go Buffs"
		end
	else if(A == 3'b111 && SW[9] == 1'b0 && KEY[1] == 1'b1)begin
		A <= 3'b000;
		counter_Enable <= 0;
		downCounter_Enable <=0;
		//downCount_Complete <=0;
		//Display High Score
		end
	else if(A == 3'b001 && downCount_Boolean == 0)begin
		downCounter_Enable <= 1'b1;
		A <= 3'b010;
		downCount_Value = LFSR_Value;
		end
	else if(A == 3'b010 && downCount_Complete == 1)begin
		counter_Enable <= 1;
		downCount_Boolean <= 0;
		downCounter_Enable <=0;
		A <= 3'b011;
		end
	else if(A == 3'b011 && KEY[1] == 1'b0)begin
		counter_Enable <= 0;
		downCounter_Enable <=0;
		//A <= 3'b100;
		//begin	
			//if({BCD3,BCD2,BCD1,BCD0} < highScore)
			//highScore <= {BCD3,BCD2,BCD1,BCD0};
		//end
		end
	//else if(A == 3'b100 && KEY[1] == 1'b0)begin
		//counter_Enable <= 0;
		//downCounter_Enable <=0;
		//A <= 3'b000;
		//end
	
	/*else begin
		//default
		A = 2'b00;
		counter_Enable = 0;
		downCounter_Enable = 0;
		downCount_Boolean = 0;
		end
	*/	
end		
		
/*	
always@(KEY[0])begin
	if(KEY[1]==0)
		ENABLE = !ENABLE;
		
	if(KEY[0]==0)
		highScore <= 0;
		A<=3'b000;
		counter_Enable <= 0;
		downCounter_Enable <= 0;
		downCount_Boolean <= 0;
		A <= 0;
end
*/

//Instantiates an instance of SevenSegment.v
//This is the decoder which translates BCD values into binary values that light the correct segments in the 7-segment display
BCD_decoder decoder_INST1(BCD0[3:0], BCD1[3:0], BCD2[3:0], BCD3[3:0], HEX0[6:0], HEX1[6:0], HEX2[6:0], HEX3[6:0]);

//Instantiates an instance of BCD_counter.v
//This code generates the values which generate numbers 1-9 for the seven-segment displays
BCD_counter BCD_Count_INST1(divided_Clock, RESET, counter_Enable, BCD3, BCD2, BCD1, BCD0);

//Instantiates an instance of Clock_divider
//This clock divides the native 50MHz clock by 25,000 to yield a 2kHz clock
clock_Divider clk_Div_INST1(MAX10_CLK1_50, divided_Clock);

//Instantiates an instance of Slow_Clock
//This clock divides the native 50MHz clock by 50,000,000 to yield a 1Hz clock
Slow_Clock Slow_Clock_INST1(MAX10_CLK1_50, Slow_Clock);

//Instantiates an instance  of LFSR 
//Generates pseudo random numbers to set the delay between pressing the start button, and the start of the timer/start indicator light
LFSR LFSR_INST1(Slow_Clock, LFSR_Value);

//instantiates an instance of down_Counter
down_Counter down_Counter_INST1(Slow_Clock, LFSR_Value, RESET, downCounter_Enable, count, downCount_Complete);
//down_Counter down_Counter_INST1(Slow_Clock, 8'b00000011, RESET, ENABLE, count, downCount_Complete);


endmodule
