//Gabriel Altman
//ECEN2350 Digital Logic
//April, 2018

//module display_MUX();